`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/05/28 14:06:23
// Design Name: 
// Module Name: MULTU
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MULTU(
 input clk,
   input [31:0]a,
   input [31:0]b,
   output reg[63:0]z
   );
  always@(*) begin
   z = (a[0] ? {32'b0,b}:64'b0)+(a[1] ? {31'b0,b,1'b0} : 64'b0)+(a[2] ? {30'b0, b, 2'b0} : 64'b0)+(a[3] ? {29'b0,b,3'b0} : 64'b0)+(a[4] ? {28'b0, b, 4'b0} : 64'b0)+(a[5] ? {27'b0,b,5'b0} : 64'b0)+(a[6] ? {26'b0, b, 6'b0} : 64'b0)+(a[7] ? {25'b0,b,7'b0} : 64'b0)+(a[8] ? {24'b0, b, 8'b0} : 64'b0)+(a[9] ? {23'b0,b,9'b0} : 64'b0)+(a[10] ? {22'b0, b, 10'b0} : 64'b0)+(a[11] ? {21'b0,b,11'b0} : 64'b0)+(a[12] ? {20'b0, b, 12'b0} : 64'b0)+(a[13] ? {19'b0,b,13'b0} : 64'b0)+(a[14] ? {18'b0, b, 14'b0} : 64'b0)+(a[15] ? {17'b0,b,15'b0} : 64'b0)+(a[16] ? {16'b0, b, 16'b0} : 64'b0)+(a[17] ? {15'b0,b,17'b0} : 64'b0)+(a[18] ? {14'b0, b, 18'b0} : 64'b0)+(a[19] ? {13'b0,b,19'b0} : 64'b0)+(a[20] ? {12'b0, b, 20'b0} : 64'b0)+(a[21] ? {11'b0,b,21'b0} : 64'b0)+(a[22] ? {10'b0, b, 22'b0} : 64'b0)+(a[23] ? {9'b0,b,23'b0} : 64'b0)+(a[24] ? {8'b0, b, 24'b0} : 64'b0)+(a[25] ? {7'b0,b,25'b0} : 64'b0)+(a[26] ? {6'b0, b, 26'b0} : 64'b0)+(a[27] ? {5'b0,b,27'b0} : 64'b0)+(a[28] ? {4'b0, b, 28'b0} : 64'b0)+(a[29] ? {3'b0,b,29'b0} : 64'b0)+(a[30] ? {2'b0, b, 30'b0} : 64'b0)+(a[31] ? {1'b0,b,31'b0} : 64'b0);
  end
endmodule
